// top_defines_fifo.sv
// Top level constant defines for fifo module
// Nosherwan Ahmed
// 17 November 2019

`define FIFO_DATA_WIDTH = 32;
`define FIFO_DEPTH = 16; 